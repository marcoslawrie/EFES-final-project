library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity testbench is
end entity;

architecture struct of testbench is


type input_DATA is array (0 to 515)
        of std_logic_vector(5 downto 0);
  constant waveform : input_DATA :=
            (           "010100",
"010111",
"100000",
"100111",
"100110",
"011110",
"010111",
"010111",
"100000",
"101000",
"101000",
"100001",
"011001",
"011000",
"011111",
"101000",
"101011",
"100101",
"011101",
"011001",
"011110",
"101000",
"101101",
"101001",
"100000",
"011011",
"011110",
"100111",
"101110",
"101100",
"100100",
"011101",
"011110",
"100110",
"101110",
"101111",
"101000",
"100000",
"011111",
"100101",
"101110",
"110001",
"101100",
"100011",
"100000",
"100101",
"101110",
"110011",
"101111",
"100111",
"100001",
"100100",
"101101",
"110100",
"110011",
"101010",
"100011",
"100100",
"101100",
"110100",
"110101",
"101110",
"100110",
"100100",
"101011",
"110100",
"110111",
"110010",
"101001",
"100101",
"101010",
"110011",
"111000",
"110101",
"101100",
"100111",
"101010",
"110010",
"111001",
"111000",
"101111",
"101000",
"101001",
"110001",
"111001",
"111010",
"110011",
"101011",
"101001",
"110000",
"111000",
"111011",
"110110",
"101101",
"101001",
"101110",
"110111",
"111100",
"111001",
"110000",
"101010",
"101101",
"110110",
"111101",
"111011",
"110011",
"101100",
"101100",
"110100",
"111100",
"111101",
"110110",
"101101",
"101100",
"110010",
"111011",
"111110",
"111000",
"101111",
"101100",
"110000",
"111001",
"111110",
"111010",
"110010",
"101100",
"101111",
"110111",
"111110",
"111100",
"110100",
"101101",
"101101",
"110101",
"111101",
"111110",
"110110",
"101110",
"101100",
"110011",
"111011",
"111110",
"111000",
"110000",
"101100",
"110000",
"111001",
"111110",
"111010",
"110001",
"101100",
"101110",
"110111",
"111101",
"111100",
"110011",
"101100",
"101100",
"110100",
"111100",
"111100",
"110101",
"101101",
"101011",
"110001",
"111010",
"111100",
"110111",
"101110",
"101010",
"101110",
"110111",
"111100",
"111000",
"101111",
"101001",
"101100",
"110100",
"111011",
"111001",
"110000",
"101001",
"101001",
"110001",
"111001",
"111001",
"110010",
"101001",
"100111",
"101110",
"110110",
"111001",
"110011",
"101010",
"100110",
"101010",
"110011",
"111000",
"110100",
"101011",
"100101",
"100111",
"110000",
"110110",
"110100",
"101100",
"100100",
"100101",
"101100",
"110100",
"110100",
"101101",
"100100",
"100010",
"101001",
"110001",
"110100",
"101110",
"100100",
"100000",
"100101",
"101110",
"110010",
"101110",
"100101",
"011111",
"100010",
"101010",
"110000",
"101110",
"100110",
"011110",
"011111",
"100110",
"101110",
"101110",
"100111",
"011110",
"011100",
"100010",
"101011",
"101101",
"100111",
"011110",
"011010",
"011111",
"100111",
"101100",
"101000",
"011111",
"011001",
"011011",
"100011",
"101010",
"101000",
"011111",
"011000",
"011000",
"100000",
"100111",
"100111",
"100000",
"010111",
"010101",
"011100",
"100100",
"100110",
"100000",
"010111",
"010011",
"011000",
"100000",
"100101",
"100001",
"011000",
"010010",
"010100",
"011101",
"100011",
"100001",
"011000",
"010001",
"010001",
"011001",
"100000",
"100001",
"011001",
"010001",
"001111",
"010101",
"011101",
"100000",
"011010",
"010001",
"001101",
"010001",
"011010",
"011111",
"011011",
"010001",
"001011",
"001110",
"010110",
"011101",
"011011",
"010010",
"001011",
"001011",
"010011",
"011010",
"011011",
"010011",
"001011",
"001001",
"001111",
"011000",
"011010",
"010100",
"001011",
"000111",
"001100",
"010101",
"011001",
"010101",
"001100",
"000110",
"001001",
"010001",
"011000",
"010110",
"001101",
"000110",
"000110",
"001110",
"010110",
"010110",
"001111",
"000110",
"000100",
"001011",
"010011",
"010110",
"010000",
"000111",
"000011",
"001000",
"010001",
"010101",
"010001",
"001000",
"000011",
"000101",
"001110",
"010100",
"010010",
"001010",
"000011",
"000011",
"001011",
"010011",
"010011",
"001100",
"000011",
"000010",
"001000",
"010001",
"010011",
"001110",
"000101",
"000001",
"000110",
"001111",
"010011",
"001111",
"000111",
"000001",
"000100",
"001100",
"010011",
"010001",
"001001",
"000001",
"000010",
"001010",
"010010",
"010010",
"001011",
"000011",
"000001",
"001000",
"010000",
"010011",
"001101",
"000101",
"000001",
"000110",
"001111",
"010011",
"010000",
"000111",
"000001",
"000100",
"001101",
"010011",
"010010",
"001001",
"000010",
"000011",
"001011",
"010011",
"010011",
"001100",
"000100",
"000010",
"001001",
"010010",
"010101",
"001111",
"000110",
"000011",
"001000",
"010001",
"010110",
"010010",
"001001",
"000100",
"000111",
"001111",
"010110",
"010100",
"001100",
"000101",
"000110",
"001110",
"010110",
"010111",
"010000",
"000111",
"000110",
"001101",
"010101",
"011000",
"010011",
"001010",
"000111",
"001100",
"010101",
"011010",
"010110",
"001101",
"001000",
"001011",
"010100",
"011011",
"011001",
"010001",
"001010",
"001011",
"010011",
"011011",
"011100",
"010101",
"001100",
"001011",
"010010",
"011011",
"011110",
"011000",
"010000",
"001100",
"010001",
"011010",
"011111",
"011100",
"010011",
"001110",
"010001",
"011010",
"100000",
"011111",
"010111",
"010000",
"010001",
"011001",
"100001",
"100010",
"011011",
"010011",
"010001",
"011000",
"100001",
"100100",
"011111",
"010110",
"010010",
"010111",
"100001",
"100110",
"100010",
"011010",
"010100",
"010111",
"100000",
"100111",
"100110",
"011110",
"010111",
"010111",
"100000",
"101000",
"101000",
"100001",
"011001",
"011000",
"011111",
"101000"
	 );
COMPONENT fir IS
	   generic (
      N_BITS_INPUT: integer := 6;
		N_BITS_COEF: integer:= 9;
		N_TAPS: integer := 17
		);
    PORT
    (
		CLK        : in  std_logic;
		RST       : in  std_logic;
		ORDER_SEL	 : in  std_logic;
		-- data input
		DATA_IN       : in  std_logic_vector( N_BITS_INPUT-1 downto 0);
		-- filtered data 
		DATA_OUT       : out std_logic_vector( N_BITS_INPUT-1 downto 0)
    );
END COMPONENT;

CONSTANT clk_period: TIME:=5 ms;

signal data_in:std_logic_vector(5 downto 0);
signal data_out:std_logic_vector( 5 downto 0);
signal CLK_TB,AUXCLK,RST_TB,ORDER_SEL_TB:std_logic;

begin

DUT: fir PORT MAP(clk_tb,rst_tb,ORDER_SEL_TB,data_in,data_out);

ClkProcess:PROCESS
BEGIN
    clk_tb<='0';
    wait for clk_period/2;
    clk_tb<='1';
    wait for clk_period/2;
END PROCESS ClkProcess;
AUXClkProcess:PROCESS
BEGIN
    AUXClk<='0';
    wait until rising_edge(clk_tb);
    AUXClk<='1';
    wait until rising_edge(clk_tb);
END PROCESS AUXClkProcess;
testProcess: PROCESS 
variable index : integer := 0;
BEGIN
data_in<="000000";
rst_tb<='0';
ORDER_SEL_TB<='1';
wait for 20 ns;
rst_tb<='1';
for k in 0 to waveform'length-1 loop
	wait until falling_edge(clk_tb);
	data_in<=waveform(index);
	index := index + 1;
end loop;



WAIT;
END PROCESS testProcess;



end architecture struct;