library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity testbench is
end entity;

architecture struct of testbench is


type input_DATA is array (0 to 507)
        of std_logic_vector(5 downto 0);
  constant waveform : input_DATA :=
            (         "100010",
    "011110",
    "011011",
    "011011",
    "100000",
    "100100",
    "100100",
    "100001",
    "011101",
    "011101",
    "100000",
    "100101",
    "100111",
    "100100",
    "100000",
    "011110",
    "100001",
    "100110",
    "101001",
    "100111",
    "100011",
    "100001",
    "100010",
    "100111",
    "101010",
    "101010",
    "100110",
    "100011",
    "100011",
    "101000",
    "101100",
    "101100",
    "101001",
    "100101",
    "100101",
    "101000",
    "101101",
    "101111",
    "101100",
    "101000",
    "100110",
    "101001",
    "101110",
    "110001",
    "101111",
    "101011",
    "101000",
    "101010",
    "101110",
    "110010",
    "110001",
    "101110",
    "101010",
    "101011",
    "101111",
    "110011",
    "110100",
    "110000",
    "101100",
    "101100",
    "101111",
    "110100",
    "110110",
    "110011",
    "101111",
    "101101",
    "110000",
    "110100",
    "110111",
    "110101",
    "110001",
    "101111",
    "110000",
    "110101",
    "111000",
    "111000",
    "110100",
    "110000",
    "110001",
    "110101",
    "111001",
    "111001",
    "110110",
    "110010",
    "110001",
    "110101",
    "111001",
    "111011",
    "111000",
    "110100",
    "110010",
    "110101",
    "111001",
    "111100",
    "111010",
    "110110",
    "110011",
    "110101",
    "111001",
    "111100",
    "111100",
    "111000",
    "110100",
    "110101",
    "111001",
    "111101",
    "111101",
    "111001",
    "110101",
    "110101",
    "111000",
    "111100",
    "111110",
    "111011",
    "110111",
    "110101",
    "110111",
    "111100",
    "111110",
    "111100",
    "111000",
    "110101",
    "110111",
    "111011",
    "111110",
    "111101",
    "111001",
    "110110",
    "110110",
    "111010",
    "111110",
    "111110",
    "111010",
    "110110",
    "110101",
    "111001",
    "111101",
    "111110",
    "111011",
    "110111",
    "110101",
    "110111",
    "111100",
    "111110",
    "111100",
    "111000",
    "110101",
    "110110",
    "111010",
    "111101",
    "111101",
    "111000",
    "110101",
    "110101",
    "111001",
    "111100",
    "111101",
    "111001",
    "110101",
    "110100",
    "110111",
    "111011",
    "111100",
    "111001",
    "110101",
    "110011",
    "110101",
    "111001",
    "111011",
    "111001",
    "110101",
    "110010",
    "110011",
    "110111",
    "111010",
    "111001",
    "110101",
    "110001",
    "110001",
    "110101",
    "111001",
    "111001",
    "110101",
    "110000",
    "101111",
    "110010",
    "110111",
    "111000",
    "110101",
    "110000",
    "101110",
    "110000",
    "110100",
    "110110",
    "110100",
    "110000",
    "101100",
    "101110",
    "110010",
    "110101",
    "110100",
    "101111",
    "101011",
    "101011",
    "101111",
    "110011",
    "110011",
    "101111",
    "101010",
    "101001",
    "101100",
    "110000",
    "110001",
    "101110",
    "101001",
    "100111",
    "101001",
    "101110",
    "110000",
    "101101",
    "101001",
    "100110",
    "100111",
    "101011",
    "101110",
    "101100",
    "101000",
    "100100",
    "100100",
    "101000",
    "101011",
    "101011",
    "100111",
    "100011",
    "100010",
    "100101",
    "101001",
    "101010",
    "100110",
    "100010",
    "011111",
    "100010",
    "100110",
    "101000",
    "100110",
    "100001",
    "011110",
    "011111",
    "100011",
    "100110",
    "100100",
    "100000",
    "011100",
    "011100",
    "100000",
    "100011",
    "100011",
    "011111",
    "011011",
    "011001",
    "011100",
    "100000",
    "100001",
    "011110",
    "011001",
    "010111",
    "011001",
    "011101",
    "100000",
    "011101",
    "011001",
    "010101",
    "010110",
    "011010",
    "011101",
    "011100",
    "011000",
    "010100",
    "010100",
    "010111",
    "011011",
    "011011",
    "010111",
    "010011",
    "010001",
    "010100",
    "011000",
    "011001",
    "010110",
    "010010",
    "001111",
    "010001",
    "010110",
    "011000",
    "010110",
    "010001",
    "001110",
    "001111",
    "010011",
    "010110",
    "010101",
    "010000",
    "001100",
    "001100",
    "010000",
    "010100",
    "010100",
    "010000",
    "001011",
    "001010",
    "001101",
    "010001",
    "010011",
    "001111",
    "001011",
    "001001",
    "001011",
    "001111",
    "010001",
    "001111",
    "001010",
    "000111",
    "001000",
    "001101",
    "010000",
    "001111",
    "001010",
    "000110",
    "000110",
    "001010",
    "001110",
    "001110",
    "001010",
    "000110",
    "000101",
    "001000",
    "001100",
    "001101",
    "001010",
    "000110",
    "000100",
    "000110",
    "001010",
    "001100",
    "001010",
    "000110",
    "000011",
    "000100",
    "001000",
    "001011",
    "001010",
    "000110",
    "000010",
    "000011",
    "000110",
    "001010",
    "001010",
    "000111",
    "000010",
    "000010",
    "000101",
    "001001",
    "001010",
    "000111",
    "000011",
    "000001",
    "000011",
    "001000",
    "001010",
    "001000",
    "000100",
    "000001",
    "000010",
    "000110",
    "001010",
    "001001",
    "000101",
    "000001",
    "000001",
    "000101",
    "001001",
    "001001",
    "000110",
    "000010",
    "000001",
    "000100",
    "001000",
    "001010",
    "000111",
    "000011",
    "000001",
    "000011",
    "001000",
    "001010",
    "001000",
    "000100",
    "000001",
    "000011",
    "000111",
    "001010",
    "001010",
    "000110",
    "000010",
    "000010",
    "000110",
    "001010",
    "001011",
    "000111",
    "000011",
    "000011",
    "000110",
    "001010",
    "001100",
    "001001",
    "000101",
    "000011",
    "000110",
    "001010",
    "001101",
    "001011",
    "000111",
    "000100",
    "000110",
    "001010",
    "001110",
    "001101",
    "001001",
    "000110",
    "000110",
    "001010",
    "001110",
    "001111",
    "001011",
    "000111",
    "000111",
    "001010",
    "001111",
    "010000",
    "001110",
    "001010",
    "001000",
    "001011",
    "001111",
    "010010",
    "010000",
    "001100",
    "001001",
    "001011",
    "010000",
    "010011",
    "010011",
    "001111",
    "001011",
    "001100",
    "010000",
    "010100",
    "010101",
    "010001",
    "001110",
    "001101",
    "010001",
    "010101",
    "010111",
    "010100",
    "010000",
    "001110",
    "010001",
    "010110",
    "011001",
    "010111",
    "010011",
    "010000",
    "010010",
    "010111",
    "011010",
    "011010",
    "010110",
    "010011",
    "010011",
    "010111",
    "011100",
    "011100",
    "011001",
    "010101",
    "010101",
    "011000",
    "011101",
    "011110",
    "011100",
    "011000",
    "010110",
    "011001",
    "011110",
    "100001",
    "011111",
    "011011",
    "011000",
    "011010",
    "011111",
    "100010",
	 "100010",
    "011110",
    "011011",
    "011011",
    "100000",
    "100100",
    "100100",
    "100001");
COMPONENT fir IS
    PORT
    (
		i_clk        : in  std_logic;
		i_rstb       : in  std_logic;
    	  -- data input
		i_data       : in  std_logic_vector( 5 downto 0);
  -- filtered data 
		o_data       : out std_logic_vector( 5 downto 0)
    );
END COMPONENT;

CONSTANT clk_period: TIME:=5 ms;

signal data_in:std_logic_vector(5 downto 0);
signal data_out:std_logic_vector( 5 downto 0);
signal clk_tb,AUXClk,rst_tb:std_logic;

begin

DUT: fir PORT MAP(clk_tb,rst_tb,data_in,data_out);

ClkProcess:PROCESS
BEGIN
    clk_tb<='0';
    wait for clk_period/2;
    clk_tb<='1';
    wait for clk_period/2;
END PROCESS ClkProcess;
AUXClkProcess:PROCESS
BEGIN
    AUXClk<='0';
    wait until rising_edge(clk_tb);
    AUXClk<='1';
    wait until rising_edge(clk_tb);
END PROCESS AUXClkProcess;
testProcess: PROCESS 
variable index : integer := 0;
BEGIN
data_in<="000000";
rst_tb<='0';
wait for 20 ns;
rst_tb<='1';
for k in 0 to waveform'length-1 loop
	wait until falling_edge(clk_tb);
	data_in<=waveform(index);
	index := index + 1;
end loop;
--wait until rising_edge(clk_tb);
--data_in<=waveform(index);
--index := index + 1;
--wait until rising_edge(clk_tb);
--data_in<=waveform(index);
--index := index + 1;
--wait until rising_edge(clk_tb);
--data_in<=waveform(index);
--index := index + 1;
--wait until rising_edge(clk_tb);
--data_in<=waveform(index);
--index := index + 1;
--wait until rising_edge(clk_tb);
--data_in<=waveform(index);
--index := index + 1;
--wait until rising_edge(clk_tb);
--data_in<=waveform(index);
--index := index + 1;
--wait until rising_edge(clk_tb);
--data_in<=waveform(index);
--index := index + 1;
--wait until rising_edge(clk_tb);
--data_in<=waveform(index);
--index := index + 1;
--wait until rising_edge(clk_tb);
--data_in<=waveform(index);
--index := index + 1;
--wait until rising_edge(clk_tb);
--data_in<=waveform(index);
--index := index + 1;



WAIT;
END PROCESS testProcess;



end architecture struct;